Library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package common_pkg is
  type std_logic_array is array (natural range <>) of std_logic_vector;
end common_pkg;
